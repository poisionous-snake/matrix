module ExpUnitFixPoint(
  input        clock,
  input        reset,
  input  [5:0] io_in_value,
  output [5:0] io_out_exp
);
  wire [5:0] x = io_in_value; // @[exp_unit.scala 81:26]
  wire [9:0] _y_T = {io_in_value, 4'h0}; // @[exp_unit.scala 82:11]
  wire [8:0] _y_T_1 = {io_in_value, 3'h0}; // @[exp_unit.scala 82:32]
  wire [9:0] _GEN_64 = {{1'd0}, _y_T_1}; // @[exp_unit.scala 82:27]
  wire [9:0] _y_T_3 = _y_T + _GEN_64; // @[exp_unit.scala 82:27]
  wire [9:0] _GEN_65 = {{4'd0}, x}; // @[exp_unit.scala 82:54]
  wire [9:0] y = _y_T_3 - _GEN_65; // @[exp_unit.scala 82:54]
  wire [7:0] v_lo = y[7:0]; // @[exp_unit.scala 85:41]
  wire [9:0] v = {2'h0,v_lo}; // @[exp_unit.scala 86:18]
  wire [9:0] _v_bits_T = {2'h0,v_lo}; // @[exp_unit.scala 62:23]
  wire [5:0] v_bits = _v_bits_T[7:2]; // @[exp_unit.scala 62:25]
  wire [9:0] _GEN_1 = v_bits == 6'h3e ? $signed(10'shfd) : $signed(10'shfe); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_2 = v_bits == 6'h3d ? $signed(10'shfc) : $signed(_GEN_1); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_3 = v_bits == 6'h3c ? $signed(10'shfa) : $signed(_GEN_2); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_4 = v_bits == 6'h3b ? $signed(10'shf9) : $signed(_GEN_3); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_5 = v_bits == 6'h3a ? $signed(10'shf8) : $signed(_GEN_4); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_6 = v_bits == 6'h39 ? $signed(10'shf7) : $signed(_GEN_5); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_7 = v_bits == 6'h38 ? $signed(10'shf6) : $signed(_GEN_6); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_8 = v_bits == 6'h37 ? $signed(10'shf4) : $signed(_GEN_7); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_9 = v_bits == 6'h36 ? $signed(10'shf3) : $signed(_GEN_8); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_10 = v_bits == 6'h35 ? $signed(10'shf2) : $signed(_GEN_9); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_11 = v_bits == 6'h34 ? $signed(10'shf2) : $signed(_GEN_10); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_12 = v_bits == 6'h33 ? $signed(10'shf1) : $signed(_GEN_11); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_13 = v_bits == 6'h32 ? $signed(10'shf0) : $signed(_GEN_12); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_14 = v_bits == 6'h31 ? $signed(10'shef) : $signed(_GEN_13); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_15 = v_bits == 6'h30 ? $signed(10'shef) : $signed(_GEN_14); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_16 = v_bits == 6'h2f ? $signed(10'shee) : $signed(_GEN_15); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_17 = v_bits == 6'h2e ? $signed(10'shed) : $signed(_GEN_16); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_18 = v_bits == 6'h2d ? $signed(10'shed) : $signed(_GEN_17); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_19 = v_bits == 6'h2c ? $signed(10'shec) : $signed(_GEN_18); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_20 = v_bits == 6'h2b ? $signed(10'shec) : $signed(_GEN_19); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_21 = v_bits == 6'h2a ? $signed(10'sheb) : $signed(_GEN_20); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_22 = v_bits == 6'h29 ? $signed(10'sheb) : $signed(_GEN_21); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_23 = v_bits == 6'h28 ? $signed(10'sheb) : $signed(_GEN_22); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_24 = v_bits == 6'h27 ? $signed(10'sheb) : $signed(_GEN_23); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_25 = v_bits == 6'h26 ? $signed(10'shea) : $signed(_GEN_24); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_26 = v_bits == 6'h25 ? $signed(10'shea) : $signed(_GEN_25); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_27 = v_bits == 6'h24 ? $signed(10'shea) : $signed(_GEN_26); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_28 = v_bits == 6'h23 ? $signed(10'shea) : $signed(_GEN_27); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_29 = v_bits == 6'h22 ? $signed(10'shea) : $signed(_GEN_28); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_30 = v_bits == 6'h21 ? $signed(10'shea) : $signed(_GEN_29); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_31 = v_bits == 6'h20 ? $signed(10'shea) : $signed(_GEN_30); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_32 = v_bits == 6'h1f ? $signed(10'shea) : $signed(_GEN_31); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_33 = v_bits == 6'h1e ? $signed(10'shea) : $signed(_GEN_32); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_34 = v_bits == 6'h1d ? $signed(10'shea) : $signed(_GEN_33); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_35 = v_bits == 6'h1c ? $signed(10'sheb) : $signed(_GEN_34); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_36 = v_bits == 6'h1b ? $signed(10'sheb) : $signed(_GEN_35); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_37 = v_bits == 6'h1a ? $signed(10'sheb) : $signed(_GEN_36); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_38 = v_bits == 6'h19 ? $signed(10'shec) : $signed(_GEN_37); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_39 = v_bits == 6'h18 ? $signed(10'shec) : $signed(_GEN_38); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_40 = v_bits == 6'h17 ? $signed(10'shec) : $signed(_GEN_39); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_41 = v_bits == 6'h16 ? $signed(10'shed) : $signed(_GEN_40); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_42 = v_bits == 6'h15 ? $signed(10'shed) : $signed(_GEN_41); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_43 = v_bits == 6'h14 ? $signed(10'shee) : $signed(_GEN_42); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_44 = v_bits == 6'h13 ? $signed(10'shee) : $signed(_GEN_43); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_45 = v_bits == 6'h12 ? $signed(10'shef) : $signed(_GEN_44); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_46 = v_bits == 6'h11 ? $signed(10'shf0) : $signed(_GEN_45); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_47 = v_bits == 6'h10 ? $signed(10'shf0) : $signed(_GEN_46); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_48 = v_bits == 6'hf ? $signed(10'shf1) : $signed(_GEN_47); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_49 = v_bits == 6'he ? $signed(10'shf2) : $signed(_GEN_48); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_50 = v_bits == 6'hd ? $signed(10'shf3) : $signed(_GEN_49); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_51 = v_bits == 6'hc ? $signed(10'shf4) : $signed(_GEN_50); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_52 = v_bits == 6'hb ? $signed(10'shf4) : $signed(_GEN_51); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_53 = v_bits == 6'ha ? $signed(10'shf5) : $signed(_GEN_52); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_54 = v_bits == 6'h9 ? $signed(10'shf6) : $signed(_GEN_53); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_55 = v_bits == 6'h8 ? $signed(10'shf7) : $signed(_GEN_54); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_56 = v_bits == 6'h7 ? $signed(10'shf8) : $signed(_GEN_55); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_57 = v_bits == 6'h6 ? $signed(10'shf9) : $signed(_GEN_56); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_58 = v_bits == 6'h5 ? $signed(10'shfa) : $signed(_GEN_57); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_59 = v_bits == 6'h4 ? $signed(10'shfb) : $signed(_GEN_58); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_60 = v_bits == 6'h3 ? $signed(10'shfc) : $signed(_GEN_59); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_61 = v_bits == 6'h2 ? $signed(10'shfe) : $signed(_GEN_60); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] _GEN_62 = v_bits == 6'h1 ? $signed(10'shff) : $signed(_GEN_61); // @[exp_unit.scala 71:46 exp_unit.scala 72:16]
  wire [9:0] d_wire = v_bits == 6'h0 ? $signed(10'sh100) : $signed(_GEN_62); // @[exp_unit.scala 67:42 exp_unit.scala 68:14]
  wire [1:0] u = y[9:8]; // @[exp_unit.scala 84:9]
  wire [9:0] z1 = $signed(v) + $signed(d_wire); // @[exp_unit.scala 88:11]
  wire [12:0] _GEN_66 = {{3{z1[9]}},z1}; // @[exp_unit.scala 89:12]
  wire [12:0] _z2_T = $signed(_GEN_66) << u; // @[exp_unit.scala 89:12]
  wire [9:0] z2 = _z2_T[9:0]; // @[exp_unit.scala 24:16 exp_unit.scala 89:6]
  assign io_out_exp = z2[9:4]; // @[exp_unit.scala 102:14]
endmodule
